module vcount(input clk, rst, sel);

    always @ (postedge clk)
        begin
            if(!rst)begin
                
            
            end
            else begin
                pass
            end
        end
    
endmodule